library ieee;
use ieee.std_logic_1164.all;

library gtlib;

entity WordMUX16to1 is
  port(Word0 : in std_logic_vector(15 downto 0);
       Word1 : in std_logic_vector(15 downto 0);
       Word2 : in std_logic_vector(15 downto 0);
       Word3 : in std_logic_vector(15 downto 0);
       Word4 : in std_logic_vector(15 downto 0);
       Word5 : in std_logic_vector(15 downto 0);
       Word6 : in std_logic_vector(15 downto 0);
       Word7 : in std_logic_vector(15 downto 0);
       Word8 : in std_logic_vector(15 downto 0);
       Word9 : in std_logic_vector(15 downto 0);
       Word10 : in std_logic_vector(15 downto 0);
       Word11 : in std_logic_vector(15 downto 0);
       Word12 : in std_logic_vector(15 downto 0);
       Word13 : in std_logic_vector(15 downto 0);
       Word14 : in std_logic_vector(15 downto 0);
       Word15 : in std_logic_vector(15 downto 0);
       sel : in std_logic_vector(3 downto 0);
       WordOut : out std_logic_vector(15 downto 0));
end WordMUX16to1;

architecture rtl of WordMUX16to1 is
  signal b33 : std_logic_vector(3 downto 0);
  signal b65 : std_logic_vector(15 downto 0);
  signal b66 : std_logic_vector(15 downto 0);
  signal b50 : std_logic_vector(15 downto 0);
  signal b51 : std_logic_vector(15 downto 0);
  signal b52 : std_logic_vector(15 downto 0);
  signal b53 : std_logic_vector(15 downto 0);
  signal b54 : std_logic_vector(15 downto 0);
  signal b55 : std_logic_vector(15 downto 0);
  signal b56 : std_logic_vector(15 downto 0);
  signal b57 : std_logic_vector(15 downto 0);
  signal b58 : std_logic_vector(15 downto 0);
  signal b59 : std_logic_vector(15 downto 0);
  signal b60 : std_logic_vector(15 downto 0);
  signal b61 : std_logic_vector(15 downto 0);
  signal b62 : std_logic_vector(15 downto 0);
  signal b63 : std_logic_vector(15 downto 0);
  signal b64 : std_logic_vector(15 downto 0);
  signal b354 : std_logic_vector(15 downto 0);
  signal b363 : std_logic_vector(15 downto 0);
  signal b364 : std_logic_vector(15 downto 0);
  signal b365 : std_logic_vector(15 downto 0);
  signal b366 : std_logic_vector(15 downto 0);
  signal b367 : std_logic_vector(15 downto 0);
  signal b368 : std_logic_vector(15 downto 0);
  signal b369 : std_logic_vector(15 downto 0);
  signal b370 : std_logic_vector(15 downto 0);
  signal w454 : std_logic;
  signal w455 : std_logic;
  signal w456 : std_logic;
  signal w457 : std_logic;
  signal w458 : std_logic;
  signal w459 : std_logic;
  signal w460 : std_logic;
  signal w461 : std_logic;
  signal b356 : std_logic_vector(15 downto 0);
  signal b359 : std_logic_vector(15 downto 0);
  signal b357 : std_logic_vector(15 downto 0);
  signal b358 : std_logic_vector(15 downto 0);
  signal b360 : std_logic_vector(15 downto 0);
  signal b361 : std_logic_vector(15 downto 0);
  signal b362 : std_logic_vector(15 downto 0);
  signal w155 : std_logic;
  signal w156 : std_logic;
  signal w173 : std_logic;
  signal w174 : std_logic;
  signal w191 : std_logic;
  signal w192 : std_logic;
  signal w209 : std_logic;
  signal w210 : std_logic;
  signal w227 : std_logic;
  signal w228 : std_logic;
  signal w245 : std_logic;
  signal w246 : std_logic;
  signal w263 : std_logic;
  signal w264 : std_logic;
  signal w281 : std_logic;
  signal w282 : std_logic;
  signal w299 : std_logic;
  signal w300 : std_logic;
  signal w317 : std_logic;
  signal w318 : std_logic;
  signal w399 : std_logic;
  signal w400 : std_logic;
  signal w417 : std_logic;
  signal w418 : std_logic;
  signal b355 : std_logic_vector(15 downto 0);
  signal b65_0_w35 : std_logic;
  signal b65_1_w36 : std_logic;
  signal b65_2_w37 : std_logic;
  signal b65_3_w38 : std_logic;
  signal b65_4_w39 : std_logic;
  signal b65_5_w40 : std_logic;
  signal b65_6_w41 : std_logic;
  signal b65_7_w42 : std_logic;
  signal b65_8_w43 : std_logic;
  signal b65_9_w44 : std_logic;
  signal b65_10_w45 : std_logic;
  signal b65_11_w46 : std_logic;
  signal b65_12_w47 : std_logic;
  signal b65_13_w48 : std_logic;
  signal b65_14_w49 : std_logic;
  signal b65_15_w50 : std_logic;
  signal b354_3_w339 : std_logic;
  signal b363_3_w332 : std_logic;
  signal b364_3_w330 : std_logic;
  signal b365_3_w329 : std_logic;
  signal b366_3_w328 : std_logic;
  signal b367_3_w327 : std_logic;
  signal b368_3_w326 : std_logic;
  signal b369_3_w325 : std_logic;
  signal b370_3_w323 : std_logic;
  signal b354_2_w324 : std_logic;
  signal b363_2_w347 : std_logic;
  signal b364_2_w346 : std_logic;
  signal b365_2_w345 : std_logic;
  signal b366_2_w344 : std_logic;
  signal b367_2_w343 : std_logic;
  signal b368_2_w342 : std_logic;
  signal b369_2_w341 : std_logic;
  signal b370_2_w340 : std_logic;
  signal b354_1_w352 : std_logic;
  signal b363_1_w363 : std_logic;
  signal b364_1_w362 : std_logic;
  signal b365_1_w361 : std_logic;
  signal b366_1_w360 : std_logic;
  signal b367_1_w359 : std_logic;
  signal b368_1_w358 : std_logic;
  signal b369_1_w357 : std_logic;
  signal b370_1_w356 : std_logic;
  signal b354_0_w389 : std_logic;
  signal b363_0_w381 : std_logic;
  signal b364_0_w378 : std_logic;
  signal b365_0_w377 : std_logic;
  signal b366_0_w376 : std_logic;
  signal b367_0_w375 : std_logic;
  signal b368_0_w374 : std_logic;
  signal b369_0_w373 : std_logic;
  signal b370_0_w372 : std_logic;
  signal b354_7_w139 : std_logic;
  signal b356_7_w140 : std_logic;
  signal b359_7_w141 : std_logic;
  signal b357_7_w142 : std_logic;
  signal b358_7_w143 : std_logic;
  signal b360_7_w144 : std_logic;
  signal b361_7_w145 : std_logic;
  signal b362_7_w146 : std_logic;
  signal b363_7_w147 : std_logic;
  signal b364_7_w148 : std_logic;
  signal b365_7_w149 : std_logic;
  signal b366_7_w150 : std_logic;
  signal b367_7_w151 : std_logic;
  signal b368_7_w152 : std_logic;
  signal b369_7_w153 : std_logic;
  signal b370_7_w154 : std_logic;
  signal b354_6_w157 : std_logic;
  signal b356_6_w158 : std_logic;
  signal b359_6_w159 : std_logic;
  signal b357_6_w160 : std_logic;
  signal b358_6_w161 : std_logic;
  signal b360_6_w162 : std_logic;
  signal b361_6_w163 : std_logic;
  signal b362_6_w164 : std_logic;
  signal b363_6_w165 : std_logic;
  signal b364_6_w166 : std_logic;
  signal b365_6_w167 : std_logic;
  signal b366_6_w168 : std_logic;
  signal b367_6_w169 : std_logic;
  signal b368_6_w170 : std_logic;
  signal b369_6_w171 : std_logic;
  signal b370_6_w172 : std_logic;
  signal b354_5_w175 : std_logic;
  signal b356_5_w176 : std_logic;
  signal b359_5_w177 : std_logic;
  signal b357_5_w178 : std_logic;
  signal b358_5_w179 : std_logic;
  signal b360_5_w180 : std_logic;
  signal b361_5_w181 : std_logic;
  signal b362_5_w182 : std_logic;
  signal b363_5_w183 : std_logic;
  signal b364_5_w184 : std_logic;
  signal b365_5_w185 : std_logic;
  signal b366_5_w186 : std_logic;
  signal b367_5_w187 : std_logic;
  signal b368_5_w188 : std_logic;
  signal b369_5_w189 : std_logic;
  signal b370_5_w190 : std_logic;
  signal b354_4_w193 : std_logic;
  signal b356_4_w194 : std_logic;
  signal b359_4_w195 : std_logic;
  signal b357_4_w196 : std_logic;
  signal b358_4_w197 : std_logic;
  signal b360_4_w198 : std_logic;
  signal b361_4_w199 : std_logic;
  signal b362_4_w200 : std_logic;
  signal b363_4_w201 : std_logic;
  signal b364_4_w202 : std_logic;
  signal b365_4_w203 : std_logic;
  signal b366_4_w204 : std_logic;
  signal b367_4_w205 : std_logic;
  signal b368_4_w206 : std_logic;
  signal b369_4_w207 : std_logic;
  signal b370_4_w208 : std_logic;
  signal b354_11_w211 : std_logic;
  signal b356_11_w212 : std_logic;
  signal b359_11_w213 : std_logic;
  signal b357_11_w214 : std_logic;
  signal b358_11_w215 : std_logic;
  signal b360_11_w216 : std_logic;
  signal b361_11_w217 : std_logic;
  signal b362_11_w218 : std_logic;
  signal b363_11_w219 : std_logic;
  signal b364_11_w220 : std_logic;
  signal b365_11_w221 : std_logic;
  signal b366_11_w222 : std_logic;
  signal b367_11_w223 : std_logic;
  signal b368_11_w224 : std_logic;
  signal b369_11_w225 : std_logic;
  signal b370_11_w226 : std_logic;
  signal b354_10_w229 : std_logic;
  signal b356_10_w230 : std_logic;
  signal b359_10_w231 : std_logic;
  signal b357_10_w232 : std_logic;
  signal b358_10_w233 : std_logic;
  signal b360_10_w234 : std_logic;
  signal b361_10_w235 : std_logic;
  signal b362_10_w236 : std_logic;
  signal b363_10_w237 : std_logic;
  signal b364_10_w238 : std_logic;
  signal b365_10_w239 : std_logic;
  signal b366_10_w240 : std_logic;
  signal b367_10_w241 : std_logic;
  signal b368_10_w242 : std_logic;
  signal b369_10_w243 : std_logic;
  signal b370_10_w244 : std_logic;
  signal b354_9_w247 : std_logic;
  signal b356_9_w248 : std_logic;
  signal b359_9_w249 : std_logic;
  signal b357_9_w250 : std_logic;
  signal b358_9_w251 : std_logic;
  signal b360_9_w252 : std_logic;
  signal b361_9_w253 : std_logic;
  signal b362_9_w254 : std_logic;
  signal b363_9_w255 : std_logic;
  signal b364_9_w256 : std_logic;
  signal b365_9_w257 : std_logic;
  signal b366_9_w258 : std_logic;
  signal b367_9_w259 : std_logic;
  signal b368_9_w260 : std_logic;
  signal b369_9_w261 : std_logic;
  signal b370_9_w262 : std_logic;
  signal b354_8_w265 : std_logic;
  signal b356_8_w266 : std_logic;
  signal b359_8_w267 : std_logic;
  signal b357_8_w268 : std_logic;
  signal b358_8_w269 : std_logic;
  signal b360_8_w270 : std_logic;
  signal b361_8_w271 : std_logic;
  signal b362_8_w272 : std_logic;
  signal b363_8_w273 : std_logic;
  signal b364_8_w274 : std_logic;
  signal b365_8_w275 : std_logic;
  signal b366_8_w276 : std_logic;
  signal b367_8_w277 : std_logic;
  signal b368_8_w278 : std_logic;
  signal b369_8_w279 : std_logic;
  signal b370_8_w280 : std_logic;
  signal b354_15_w283 : std_logic;
  signal b356_15_w284 : std_logic;
  signal b359_15_w285 : std_logic;
  signal b357_15_w286 : std_logic;
  signal b358_15_w287 : std_logic;
  signal b360_15_w288 : std_logic;
  signal b361_15_w289 : std_logic;
  signal b362_15_w290 : std_logic;
  signal b363_15_w291 : std_logic;
  signal b364_15_w292 : std_logic;
  signal b365_15_w293 : std_logic;
  signal b366_15_w294 : std_logic;
  signal b367_15_w295 : std_logic;
  signal b368_15_w296 : std_logic;
  signal b369_15_w297 : std_logic;
  signal b370_15_w298 : std_logic;
  signal b354_14_w301 : std_logic;
  signal b356_14_w302 : std_logic;
  signal b359_14_w303 : std_logic;
  signal b357_14_w304 : std_logic;
  signal b358_14_w305 : std_logic;
  signal b360_14_w306 : std_logic;
  signal b361_14_w307 : std_logic;
  signal b362_14_w308 : std_logic;
  signal b363_14_w309 : std_logic;
  signal b364_14_w310 : std_logic;
  signal b365_14_w311 : std_logic;
  signal b366_14_w312 : std_logic;
  signal b367_14_w313 : std_logic;
  signal b368_14_w314 : std_logic;
  signal b369_14_w315 : std_logic;
  signal b370_14_w316 : std_logic;
  signal b354_13_w319 : std_logic;
  signal b356_13_w320 : std_logic;
  signal b359_13_w321 : std_logic;
  signal b357_13_w322 : std_logic;
  signal b358_13_w368 : std_logic;
  signal b360_13_w379 : std_logic;
  signal b361_13_w380 : std_logic;
  signal b362_13_w390 : std_logic;
  signal b363_13_w391 : std_logic;
  signal b364_13_w392 : std_logic;
  signal b365_13_w393 : std_logic;
  signal b366_13_w394 : std_logic;
  signal b367_13_w395 : std_logic;
  signal b368_13_w396 : std_logic;
  signal b369_13_w397 : std_logic;
  signal b370_13_w398 : std_logic;
  signal b354_12_w401 : std_logic;
  signal b356_12_w402 : std_logic;
  signal b359_12_w403 : std_logic;
  signal b357_12_w404 : std_logic;
  signal b358_12_w405 : std_logic;
  signal b360_12_w406 : std_logic;
  signal b361_12_w407 : std_logic;
  signal b362_12_w408 : std_logic;
  signal b363_12_w409 : std_logic;
  signal b364_12_w410 : std_logic;
  signal b365_12_w411 : std_logic;
  signal b366_12_w412 : std_logic;
  signal b367_12_w413 : std_logic;
  signal b368_12_w414 : std_logic;
  signal b369_12_w415 : std_logic;
  signal b370_12_w416 : std_logic;
  signal b355_0 : std_logic;
  signal b355_1 : std_logic;
  signal b355_2 : std_logic;
  signal b355_3 : std_logic;
  signal b355_4 : std_logic;
  signal b355_5 : std_logic;
  signal b355_6 : std_logic;
  signal b355_7 : std_logic;
  signal b355_8 : std_logic;
  signal b355_9 : std_logic;
  signal b355_10 : std_logic;
  signal b355_11 : std_logic;
  signal b355_12 : std_logic;
  signal b355_13 : std_logic;
  signal b355_14 : std_logic;
  signal b356_0_w388 : std_logic;
  signal b359_0_w387 : std_logic;
  signal b357_0_w386 : std_logic;
  signal b358_0_w385 : std_logic;
  signal b360_0_w384 : std_logic;
  signal b361_0_w383 : std_logic;
  signal b362_0_w382 : std_logic;
  signal b356_1_w371 : std_logic;
  signal b359_1_w370 : std_logic;
  signal b357_1_w369 : std_logic;
  signal b358_1_w367 : std_logic;
  signal b360_1_w366 : std_logic;
  signal b361_1_w365 : std_logic;
  signal b362_1_w364 : std_logic;
  signal b356_2_w355 : std_logic;
  signal b359_2_w436 : std_logic;
  signal b357_2_w437 : std_logic;
  signal b358_2_w438 : std_logic;
  signal b360_2_w439 : std_logic;
  signal b361_2_w440 : std_logic;
  signal b362_2_w441 : std_logic;
  signal b356_3_w442 : std_logic;
  signal b359_3_w443 : std_logic;
  signal b357_3_w444 : std_logic;
  signal b358_3_w445 : std_logic;
  signal b360_3_w446 : std_logic;
  signal b361_3_w447 : std_logic;
  signal b362_3_w448 : std_logic;
  signal b355_15 : std_logic;

  component Decoder4to16
    port(DecIn : in std_logic_vector(3 downto 0);
         DecOut : out std_logic_vector(15 downto 0));
  end component;

  component GT_OR8
    port(A : in std_logic;
         B : in std_logic;
         C : in std_logic;
         D : in std_logic;
         E : in std_logic;
         F : in std_logic;
         G : in std_logic;
         H : in std_logic;
         Z : out std_logic);
  end component;

  component GT_OR2
    port(A : in std_logic;
         B : in std_logic;
         Z : out std_logic);
  end component;

  component WordSelector
    port(WordIn : in std_logic_vector(15 downto 0);
         sel : in std_logic;
         WordOut : out std_logic_vector(15 downto 0));
  end component;

begin
  b66 <= Word0;
  b50 <= Word1;
  b51 <= Word2;
  b52 <= Word3;
  b53 <= Word4;
  b54 <= Word5;
  b55 <= Word6;
  b56 <= Word7;
  b57 <= Word8;
  b58 <= Word9;
  b59 <= Word10;
  b60 <= Word11;
  b61 <= Word12;
  b62 <= Word13;
  b63 <= Word14;
  b64 <= Word15;
  b33 <= sel;
  WordOut <= b355;

  b355(15) <= b355_15;
  b355(14) <= b355_14;
  b355(13) <= b355_13;
  b355(12) <= b355_12;
  b355(11) <= b355_11;
  b355(10) <= b355_10;
  b355(9) <= b355_9;
  b355(8) <= b355_8;
  b355(7) <= b355_7;
  b355(6) <= b355_6;
  b355(5) <= b355_5;
  b355(4) <= b355_4;
  b355(3) <= b355_3;
  b355(2) <= b355_2;
  b355(1) <= b355_1;
  b355(0) <= b355_0;

  b65_0_w35 <= b65(0);
  b65_1_w36 <= b65(1);
  b65_2_w37 <= b65(2);
  b65_3_w38 <= b65(3);
  b65_4_w39 <= b65(4);
  b65_5_w40 <= b65(5);
  b65_6_w41 <= b65(6);
  b65_7_w42 <= b65(7);
  b65_8_w43 <= b65(8);
  b65_9_w44 <= b65(9);
  b65_10_w45 <= b65(10);
  b65_11_w46 <= b65(11);
  b65_12_w47 <= b65(12);
  b65_13_w48 <= b65(13);
  b65_14_w49 <= b65(14);
  b65_15_w50 <= b65(15);
  b354_3_w339 <= b354(3);
  b363_3_w332 <= b363(3);
  b364_3_w330 <= b364(3);
  b365_3_w329 <= b365(3);
  b366_3_w328 <= b366(3);
  b367_3_w327 <= b367(3);
  b368_3_w326 <= b368(3);
  b369_3_w325 <= b369(3);
  b370_3_w323 <= b370(3);
  b354_2_w324 <= b354(2);
  b363_2_w347 <= b363(2);
  b364_2_w346 <= b364(2);
  b365_2_w345 <= b365(2);
  b366_2_w344 <= b366(2);
  b367_2_w343 <= b367(2);
  b368_2_w342 <= b368(2);
  b369_2_w341 <= b369(2);
  b370_2_w340 <= b370(2);
  b354_1_w352 <= b354(1);
  b363_1_w363 <= b363(1);
  b364_1_w362 <= b364(1);
  b365_1_w361 <= b365(1);
  b366_1_w360 <= b366(1);
  b367_1_w359 <= b367(1);
  b368_1_w358 <= b368(1);
  b369_1_w357 <= b369(1);
  b370_1_w356 <= b370(1);
  b354_0_w389 <= b354(0);
  b363_0_w381 <= b363(0);
  b364_0_w378 <= b364(0);
  b365_0_w377 <= b365(0);
  b366_0_w376 <= b366(0);
  b367_0_w375 <= b367(0);
  b368_0_w374 <= b368(0);
  b369_0_w373 <= b369(0);
  b370_0_w372 <= b370(0);
  b354_7_w139 <= b354(7);
  b356_7_w140 <= b356(7);
  b359_7_w141 <= b359(7);
  b357_7_w142 <= b357(7);
  b358_7_w143 <= b358(7);
  b360_7_w144 <= b360(7);
  b361_7_w145 <= b361(7);
  b362_7_w146 <= b362(7);
  b363_7_w147 <= b363(7);
  b364_7_w148 <= b364(7);
  b365_7_w149 <= b365(7);
  b366_7_w150 <= b366(7);
  b367_7_w151 <= b367(7);
  b368_7_w152 <= b368(7);
  b369_7_w153 <= b369(7);
  b370_7_w154 <= b370(7);
  b354_6_w157 <= b354(6);
  b356_6_w158 <= b356(6);
  b359_6_w159 <= b359(6);
  b357_6_w160 <= b357(6);
  b358_6_w161 <= b358(6);
  b360_6_w162 <= b360(6);
  b361_6_w163 <= b361(6);
  b362_6_w164 <= b362(6);
  b363_6_w165 <= b363(6);
  b364_6_w166 <= b364(6);
  b365_6_w167 <= b365(6);
  b366_6_w168 <= b366(6);
  b367_6_w169 <= b367(6);
  b368_6_w170 <= b368(6);
  b369_6_w171 <= b369(6);
  b370_6_w172 <= b370(6);
  b354_5_w175 <= b354(5);
  b356_5_w176 <= b356(5);
  b359_5_w177 <= b359(5);
  b357_5_w178 <= b357(5);
  b358_5_w179 <= b358(5);
  b360_5_w180 <= b360(5);
  b361_5_w181 <= b361(5);
  b362_5_w182 <= b362(5);
  b363_5_w183 <= b363(5);
  b364_5_w184 <= b364(5);
  b365_5_w185 <= b365(5);
  b366_5_w186 <= b366(5);
  b367_5_w187 <= b367(5);
  b368_5_w188 <= b368(5);
  b369_5_w189 <= b369(5);
  b370_5_w190 <= b370(5);
  b354_4_w193 <= b354(4);
  b356_4_w194 <= b356(4);
  b359_4_w195 <= b359(4);
  b357_4_w196 <= b357(4);
  b358_4_w197 <= b358(4);
  b360_4_w198 <= b360(4);
  b361_4_w199 <= b361(4);
  b362_4_w200 <= b362(4);
  b363_4_w201 <= b363(4);
  b364_4_w202 <= b364(4);
  b365_4_w203 <= b365(4);
  b366_4_w204 <= b366(4);
  b367_4_w205 <= b367(4);
  b368_4_w206 <= b368(4);
  b369_4_w207 <= b369(4);
  b370_4_w208 <= b370(4);
  b354_11_w211 <= b354(11);
  b356_11_w212 <= b356(11);
  b359_11_w213 <= b359(11);
  b357_11_w214 <= b357(11);
  b358_11_w215 <= b358(11);
  b360_11_w216 <= b360(11);
  b361_11_w217 <= b361(11);
  b362_11_w218 <= b362(11);
  b363_11_w219 <= b363(11);
  b364_11_w220 <= b364(11);
  b365_11_w221 <= b365(11);
  b366_11_w222 <= b366(11);
  b367_11_w223 <= b367(11);
  b368_11_w224 <= b368(11);
  b369_11_w225 <= b369(11);
  b370_11_w226 <= b370(11);
  b354_10_w229 <= b354(10);
  b356_10_w230 <= b356(10);
  b359_10_w231 <= b359(10);
  b357_10_w232 <= b357(10);
  b358_10_w233 <= b358(10);
  b360_10_w234 <= b360(10);
  b361_10_w235 <= b361(10);
  b362_10_w236 <= b362(10);
  b363_10_w237 <= b363(10);
  b364_10_w238 <= b364(10);
  b365_10_w239 <= b365(10);
  b366_10_w240 <= b366(10);
  b367_10_w241 <= b367(10);
  b368_10_w242 <= b368(10);
  b369_10_w243 <= b369(10);
  b370_10_w244 <= b370(10);
  b354_9_w247 <= b354(9);
  b356_9_w248 <= b356(9);
  b359_9_w249 <= b359(9);
  b357_9_w250 <= b357(9);
  b358_9_w251 <= b358(9);
  b360_9_w252 <= b360(9);
  b361_9_w253 <= b361(9);
  b362_9_w254 <= b362(9);
  b363_9_w255 <= b363(9);
  b364_9_w256 <= b364(9);
  b365_9_w257 <= b365(9);
  b366_9_w258 <= b366(9);
  b367_9_w259 <= b367(9);
  b368_9_w260 <= b368(9);
  b369_9_w261 <= b369(9);
  b370_9_w262 <= b370(9);
  b354_8_w265 <= b354(8);
  b356_8_w266 <= b356(8);
  b359_8_w267 <= b359(8);
  b357_8_w268 <= b357(8);
  b358_8_w269 <= b358(8);
  b360_8_w270 <= b360(8);
  b361_8_w271 <= b361(8);
  b362_8_w272 <= b362(8);
  b363_8_w273 <= b363(8);
  b364_8_w274 <= b364(8);
  b365_8_w275 <= b365(8);
  b366_8_w276 <= b366(8);
  b367_8_w277 <= b367(8);
  b368_8_w278 <= b368(8);
  b369_8_w279 <= b369(8);
  b370_8_w280 <= b370(8);
  b354_15_w283 <= b354(15);
  b356_15_w284 <= b356(15);
  b359_15_w285 <= b359(15);
  b357_15_w286 <= b357(15);
  b358_15_w287 <= b358(15);
  b360_15_w288 <= b360(15);
  b361_15_w289 <= b361(15);
  b362_15_w290 <= b362(15);
  b363_15_w291 <= b363(15);
  b364_15_w292 <= b364(15);
  b365_15_w293 <= b365(15);
  b366_15_w294 <= b366(15);
  b367_15_w295 <= b367(15);
  b368_15_w296 <= b368(15);
  b369_15_w297 <= b369(15);
  b370_15_w298 <= b370(15);
  b354_14_w301 <= b354(14);
  b356_14_w302 <= b356(14);
  b359_14_w303 <= b359(14);
  b357_14_w304 <= b357(14);
  b358_14_w305 <= b358(14);
  b360_14_w306 <= b360(14);
  b361_14_w307 <= b361(14);
  b362_14_w308 <= b362(14);
  b363_14_w309 <= b363(14);
  b364_14_w310 <= b364(14);
  b365_14_w311 <= b365(14);
  b366_14_w312 <= b366(14);
  b367_14_w313 <= b367(14);
  b368_14_w314 <= b368(14);
  b369_14_w315 <= b369(14);
  b370_14_w316 <= b370(14);
  b354_13_w319 <= b354(13);
  b356_13_w320 <= b356(13);
  b359_13_w321 <= b359(13);
  b357_13_w322 <= b357(13);
  b358_13_w368 <= b358(13);
  b360_13_w379 <= b360(13);
  b361_13_w380 <= b361(13);
  b362_13_w390 <= b362(13);
  b363_13_w391 <= b363(13);
  b364_13_w392 <= b364(13);
  b365_13_w393 <= b365(13);
  b366_13_w394 <= b366(13);
  b367_13_w395 <= b367(13);
  b368_13_w396 <= b368(13);
  b369_13_w397 <= b369(13);
  b370_13_w398 <= b370(13);
  b354_12_w401 <= b354(12);
  b356_12_w402 <= b356(12);
  b359_12_w403 <= b359(12);
  b357_12_w404 <= b357(12);
  b358_12_w405 <= b358(12);
  b360_12_w406 <= b360(12);
  b361_12_w407 <= b361(12);
  b362_12_w408 <= b362(12);
  b363_12_w409 <= b363(12);
  b364_12_w410 <= b364(12);
  b365_12_w411 <= b365(12);
  b366_12_w412 <= b366(12);
  b367_12_w413 <= b367(12);
  b368_12_w414 <= b368(12);
  b369_12_w415 <= b369(12);
  b370_12_w416 <= b370(12);
  b356_0_w388 <= b356(0);
  b359_0_w387 <= b359(0);
  b357_0_w386 <= b357(0);
  b358_0_w385 <= b358(0);
  b360_0_w384 <= b360(0);
  b361_0_w383 <= b361(0);
  b362_0_w382 <= b362(0);
  b356_1_w371 <= b356(1);
  b359_1_w370 <= b359(1);
  b357_1_w369 <= b357(1);
  b358_1_w367 <= b358(1);
  b360_1_w366 <= b360(1);
  b361_1_w365 <= b361(1);
  b362_1_w364 <= b362(1);
  b356_2_w355 <= b356(2);
  b359_2_w436 <= b359(2);
  b357_2_w437 <= b357(2);
  b358_2_w438 <= b358(2);
  b360_2_w439 <= b360(2);
  b361_2_w440 <= b361(2);
  b362_2_w441 <= b362(2);
  b356_3_w442 <= b356(3);
  b359_3_w443 <= b359(3);
  b357_3_w444 <= b357(3);
  b358_3_w445 <= b358(3);
  b360_3_w446 <= b360(3);
  b361_3_w447 <= b361(3);
  b362_3_w448 <= b362(3);

  s1 : Decoder4to16
    port map(
      DecIn => b33,
      DecOut => b65);

  s19 : GT_OR8
    port map(
      A => b363_3_w332,
      B => b364_3_w330,
      C => b365_3_w329,
      D => b366_3_w328,
      E => b367_3_w327,
      F => b368_3_w326,
      G => b369_3_w325,
      H => b370_3_w323,
      Z => w455);

  s18 : GT_OR8
    port map(
      A => b354_3_w339,
      Z => w454,
      B => b356_3_w442,
      C => b359_3_w443,
      D => b357_3_w444,
      E => b358_3_w445,
      F => b360_3_w446,
      G => b361_3_w447,
      H => b362_3_w448);

  s20 : GT_OR2
    port map(
      A => w454,
      B => w455,
      Z => b355_3);

  s24 : GT_OR8
    port map(
      A => b363_1_w363,
      B => b364_1_w362,
      C => b365_1_w361,
      D => b366_1_w360,
      E => b367_1_w359,
      F => b368_1_w358,
      G => b369_1_w357,
      H => b370_1_w356,
      Z => w458);

  s25 : GT_OR8
    port map(
      A => b354_1_w352,
      Z => w459,
      B => b356_1_w371,
      C => b359_1_w370,
      D => b357_1_w369,
      E => b358_1_w367,
      F => b360_1_w366,
      G => b361_1_w365,
      H => b362_1_w364);

  s26 : GT_OR2
    port map(
      B => w458,
      A => w459,
      Z => b355_1);

  s27 : GT_OR8
    port map(
      A => b363_0_w381,
      B => b364_0_w378,
      C => b365_0_w377,
      D => b366_0_w376,
      E => b367_0_w375,
      F => b368_0_w374,
      G => b369_0_w373,
      H => b370_0_w372,
      Z => w461);

  s28 : GT_OR8
    port map(
      A => b354_0_w389,
      Z => w460,
      B => b356_0_w388,
      C => b359_0_w387,
      D => b357_0_w386,
      E => b358_0_w385,
      F => b360_0_w384,
      G => b361_0_w383,
      H => b362_0_w382);

  s29 : GT_OR2
    port map(
      A => w460,
      B => w461,
      Z => b355_0);

  s21 : GT_OR8
    port map(
      A => b363_2_w347,
      B => b364_2_w346,
      C => b365_2_w345,
      D => b366_2_w344,
      E => b367_2_w343,
      F => b368_2_w342,
      G => b369_2_w341,
      H => b370_2_w340,
      Z => w457);

  s22 : GT_OR8
    port map(
      A => b354_2_w324,
      Z => w456,
      B => b356_2_w355,
      C => b359_2_w436,
      D => b357_2_w437,
      E => b358_2_w438,
      F => b360_2_w439,
      G => b361_2_w440,
      H => b362_2_w441);

  s23 : GT_OR2
    port map(
      A => w456,
      B => w457,
      Z => b355_2);

  s30 : GT_OR8
    port map(
      A => b363_7_w147,
      B => b364_7_w148,
      C => b365_7_w149,
      D => b366_7_w150,
      E => b367_7_w151,
      F => b368_7_w152,
      G => b369_7_w153,
      H => b370_7_w154,
      Z => w156);

  s31 : GT_OR8
    port map(
      A => b354_7_w139,
      B => b356_7_w140,
      C => b359_7_w141,
      D => b357_7_w142,
      E => b358_7_w143,
      F => b360_7_w144,
      G => b361_7_w145,
      H => b362_7_w146,
      Z => w155);

  s32 : GT_OR2
    port map(
      A => w155,
      B => w156,
      Z => b355_7);

  s33 : GT_OR8
    port map(
      A => b363_5_w183,
      B => b364_5_w184,
      C => b365_5_w185,
      D => b366_5_w186,
      E => b367_5_w187,
      F => b368_5_w188,
      G => b369_5_w189,
      H => b370_5_w190,
      Z => w191);

  s34 : GT_OR8
    port map(
      A => b354_5_w175,
      B => b356_5_w176,
      C => b359_5_w177,
      D => b357_5_w178,
      E => b358_5_w179,
      F => b360_5_w180,
      G => b361_5_w181,
      H => b362_5_w182,
      Z => w192);

  s35 : GT_OR2
    port map(
      B => w191,
      A => w192,
      Z => b355_5);

  s36 : GT_OR8
    port map(
      A => b363_4_w201,
      B => b364_4_w202,
      C => b365_4_w203,
      D => b366_4_w204,
      E => b367_4_w205,
      F => b368_4_w206,
      G => b369_4_w207,
      H => b370_4_w208,
      Z => w210);

  s37 : GT_OR8
    port map(
      A => b354_4_w193,
      B => b356_4_w194,
      C => b359_4_w195,
      D => b357_4_w196,
      E => b358_4_w197,
      F => b360_4_w198,
      G => b361_4_w199,
      H => b362_4_w200,
      Z => w209);

  s38 : GT_OR2
    port map(
      A => w209,
      B => w210,
      Z => b355_4);

  s39 : GT_OR8
    port map(
      A => b363_6_w165,
      B => b364_6_w166,
      C => b365_6_w167,
      D => b366_6_w168,
      E => b367_6_w169,
      F => b368_6_w170,
      G => b369_6_w171,
      H => b370_6_w172,
      Z => w174);

  s40 : GT_OR8
    port map(
      A => b354_6_w157,
      B => b356_6_w158,
      C => b359_6_w159,
      D => b357_6_w160,
      E => b358_6_w161,
      F => b360_6_w162,
      G => b361_6_w163,
      H => b362_6_w164,
      Z => w173);

  s41 : GT_OR2
    port map(
      A => w173,
      B => w174,
      Z => b355_6);

  s42 : GT_OR8
    port map(
      A => b363_11_w219,
      B => b364_11_w220,
      C => b365_11_w221,
      D => b366_11_w222,
      E => b367_11_w223,
      F => b368_11_w224,
      G => b369_11_w225,
      H => b370_11_w226,
      Z => w228);

  s43 : GT_OR8
    port map(
      A => b354_11_w211,
      B => b356_11_w212,
      C => b359_11_w213,
      D => b357_11_w214,
      E => b358_11_w215,
      F => b360_11_w216,
      G => b361_11_w217,
      H => b362_11_w218,
      Z => w227);

  s44 : GT_OR2
    port map(
      A => w227,
      B => w228,
      Z => b355_11);

  s45 : GT_OR8
    port map(
      A => b363_9_w255,
      B => b364_9_w256,
      C => b365_9_w257,
      D => b366_9_w258,
      E => b367_9_w259,
      F => b368_9_w260,
      G => b369_9_w261,
      H => b370_9_w262,
      Z => w263);

  s46 : GT_OR8
    port map(
      A => b354_9_w247,
      B => b356_9_w248,
      C => b359_9_w249,
      D => b357_9_w250,
      E => b358_9_w251,
      F => b360_9_w252,
      G => b361_9_w253,
      H => b362_9_w254,
      Z => w264);

  s47 : GT_OR2
    port map(
      B => w263,
      A => w264,
      Z => b355_9);

  s48 : GT_OR8
    port map(
      A => b363_8_w273,
      B => b364_8_w274,
      C => b365_8_w275,
      D => b366_8_w276,
      E => b367_8_w277,
      F => b368_8_w278,
      G => b369_8_w279,
      H => b370_8_w280,
      Z => w282);

  s49 : GT_OR8
    port map(
      A => b354_8_w265,
      B => b356_8_w266,
      C => b359_8_w267,
      D => b357_8_w268,
      E => b358_8_w269,
      F => b360_8_w270,
      G => b361_8_w271,
      H => b362_8_w272,
      Z => w281);

  s50 : GT_OR2
    port map(
      A => w281,
      B => w282,
      Z => b355_8);

  s51 : GT_OR8
    port map(
      A => b363_10_w237,
      B => b364_10_w238,
      C => b365_10_w239,
      D => b366_10_w240,
      E => b367_10_w241,
      F => b368_10_w242,
      G => b369_10_w243,
      H => b370_10_w244,
      Z => w246);

  s52 : GT_OR8
    port map(
      A => b354_10_w229,
      B => b356_10_w230,
      C => b359_10_w231,
      D => b357_10_w232,
      E => b358_10_w233,
      F => b360_10_w234,
      G => b361_10_w235,
      H => b362_10_w236,
      Z => w245);

  s53 : GT_OR2
    port map(
      A => w245,
      B => w246,
      Z => b355_10);

  s54 : GT_OR8
    port map(
      A => b363_15_w291,
      B => b364_15_w292,
      C => b365_15_w293,
      D => b366_15_w294,
      E => b367_15_w295,
      F => b368_15_w296,
      G => b369_15_w297,
      H => b370_15_w298,
      Z => w300);

  s55 : GT_OR8
    port map(
      A => b354_15_w283,
      B => b356_15_w284,
      C => b359_15_w285,
      D => b357_15_w286,
      E => b358_15_w287,
      F => b360_15_w288,
      G => b361_15_w289,
      H => b362_15_w290,
      Z => w299);

  s56 : GT_OR2
    port map(
      A => w299,
      B => w300,
      Z => b355_15);

  s57 : GT_OR8
    port map(
      A => b363_13_w391,
      B => b364_13_w392,
      C => b365_13_w393,
      D => b366_13_w394,
      E => b367_13_w395,
      F => b368_13_w396,
      G => b369_13_w397,
      H => b370_13_w398,
      Z => w399);

  s58 : GT_OR8
    port map(
      A => b354_13_w319,
      B => b356_13_w320,
      C => b359_13_w321,
      D => b357_13_w322,
      E => b358_13_w368,
      F => b360_13_w379,
      G => b361_13_w380,
      H => b362_13_w390,
      Z => w400);

  s59 : GT_OR2
    port map(
      B => w399,
      A => w400,
      Z => b355_13);

  s60 : GT_OR8
    port map(
      A => b363_12_w409,
      B => b364_12_w410,
      C => b365_12_w411,
      D => b366_12_w412,
      E => b367_12_w413,
      F => b368_12_w414,
      G => b369_12_w415,
      H => b370_12_w416,
      Z => w418);

  s61 : GT_OR8
    port map(
      A => b354_12_w401,
      B => b356_12_w402,
      C => b359_12_w403,
      D => b357_12_w404,
      E => b358_12_w405,
      F => b360_12_w406,
      G => b361_12_w407,
      H => b362_12_w408,
      Z => w417);

  s62 : GT_OR2
    port map(
      A => w417,
      B => w418,
      Z => b355_12);

  s63 : GT_OR8
    port map(
      A => b363_14_w309,
      B => b364_14_w310,
      C => b365_14_w311,
      D => b366_14_w312,
      E => b367_14_w313,
      F => b368_14_w314,
      G => b369_14_w315,
      H => b370_14_w316,
      Z => w318);

  s64 : GT_OR8
    port map(
      A => b354_14_w301,
      B => b356_14_w302,
      C => b359_14_w303,
      D => b357_14_w304,
      E => b358_14_w305,
      F => b360_14_w306,
      G => b361_14_w307,
      H => b362_14_w308,
      Z => w317);

  s65 : GT_OR2
    port map(
      A => w317,
      B => w318,
      Z => b355_14);

  s66 : WordSelector
    port map(
      sel => b65_0_w35,
      WordIn => b66,
      WordOut => b370);

  s67 : WordSelector
    port map(
      sel => b65_1_w36,
      WordIn => b50,
      WordOut => b369);

  s68 : WordSelector
    port map(
      sel => b65_2_w37,
      WordIn => b51,
      WordOut => b368);

  s69 : WordSelector
    port map(
      sel => b65_3_w38,
      WordIn => b52,
      WordOut => b367);

  s70 : WordSelector
    port map(
      sel => b65_4_w39,
      WordIn => b53,
      WordOut => b366);

  s71 : WordSelector
    port map(
      sel => b65_5_w40,
      WordIn => b54,
      WordOut => b365);

  s72 : WordSelector
    port map(
      sel => b65_6_w41,
      WordIn => b55,
      WordOut => b364);

  s73 : WordSelector
    port map(
      sel => b65_7_w42,
      WordIn => b56,
      WordOut => b363);

  s74 : WordSelector
    port map(
      sel => b65_8_w43,
      WordIn => b57,
      WordOut => b362);

  s75 : WordSelector
    port map(
      sel => b65_9_w44,
      WordIn => b58,
      WordOut => b361);

  s76 : WordSelector
    port map(
      sel => b65_10_w45,
      WordIn => b59,
      WordOut => b360);

  s77 : WordSelector
    port map(
      sel => b65_11_w46,
      WordIn => b60,
      WordOut => b358);

  s78 : WordSelector
    port map(
      sel => b65_12_w47,
      WordIn => b61,
      WordOut => b357);

  s79 : WordSelector
    port map(
      sel => b65_13_w48,
      WordIn => b62,
      WordOut => b359);

  s80 : WordSelector
    port map(
      sel => b65_14_w49,
      WordIn => b63,
      WordOut => b356);

  s81 : WordSelector
    port map(
      sel => b65_15_w50,
      WordIn => b64,
      WordOut => b354);

end rtl;

